LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
USE ieee.std_logic_unsigned.all ;

entity mux_21 is
	port (Sel	: in STD_LOGIC;
		  A		: in STD_LOGIC_VECTOR (31 downto 0);
		  B		: in STD_LOGIC_VECTOR (31 downto 0);
		  X		: out STD_LOGIC_VECTOR (31 downto 0));
end mux_21;

architecture mux_21_arch of mux_21 is
begin
	X <= A when (Sel = '1') else B;
end mux_21_arch;