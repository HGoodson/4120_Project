library ieee;
use ieee.std_logic_1164.all;

package DFFout is
  type DFFArray is array (natural range <>) of std_logic_vector(31 DOWNTO 0);
end package;

package body DFFout is
end package body;
